/* 
Copyright (c) 2018, IIT Madras All rights reserved.

Redistribution and use in source and binary forms, with or without modification, are permitted
provided that the following conditions are met:

* Redistributions of source code must retain the above copyright notice, this list of conditions
  and the following disclaimer.  
* Redistributions in binary form must reproduce the above copyright notice, this list of 
  conditions and the following disclaimer in the documentation and/or other materials provided 
 with the distribution.  
* Neither the name of IIT Madras  nor the names of its contributors may be used to endorse or 
  promote products derived from this software without specific prior written permission.

THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS
OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR
CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE,
DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER
IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT 
OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
--------------------------------------------------------------------------------------------------

Author: Gokulan Ravi
Email id: gokulan97@gmail.com
Details:

--------------------------------------------------------------------------------------------------
*/

package systolic_tb;
  imoprt systolic::*;
  import unified_buffer::*;

  `include  "systolic.defines"

  interface Ifc_systolic_tb#(numeric type entry_width,
                             numeric type num_entries,
                             numeric type log_num_entries,
                             numeric type num_banks,
                             numeric type num_buffers.
                             numeric type num_rows,
                             numeric type num_cols,
                             numeric type mul_width);

  endinterface

  module mksystolic_tb(Ifc_systolic_tb#(entry_width,
                                        num_entries,
                                        log_num_entries,
                                        num_banks,
                                        num_buffers,
                                        num_rows,
                                        num_cols,
                                        mul_width));

    let numRows = valueOf(num_rows);
    let numCols = valueOf(num_cols);
    let numBuffers = valueOf(num_buffers);

    Ifc_systolic#(num_rows, num_cols, mul_width) systolic <- mksystolic;
    Ifc_unified_buffer#(entry_width, num_entries, log_num_entries, num_banks, num_buffers) buffers <- mkunified_buffer;

    for(Integer i=0; i<numRows; i=i+1)begin
      for(Integer j=0; j<numBuffers; j=j+1)begin
        rule rl_always_fire;
          let val <- buffers[j][i].get();
          rfifo[i].send_rowbuf_value(tagged Valid val);
        endrule
      end
    end


  endmodule



endpackage
